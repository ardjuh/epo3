l
2
hoi
