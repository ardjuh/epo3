library IEEE;
use IEEE.std_logic_1164.ALL;

entity main is
   port(        clk    : in  std_logic;
        reset  : in  std_logic;
        vga_hsync : out std_logic;
        vga_vsync : out std_logic;
        r   : out std_logic_vector(3 downto 0);
        g : out std_logic_vector(3 downto 0);
        b  : out std_logic_vector(3 downto 0);
	screentype : in std_logic_vector (1 downto 0);
	cursor : in std_logic_vector (2 downto 0);
	
	player	: in std_logic_vector (2 downto 0);

	player_a : in std_logic;
        card1_1 : in std_logic_vector (3 downto 0);
        card1_2 : in std_logic_vector (3 downto 0);
        card1_3 : in std_logic_vector (3 downto 0);
        card1_4 : in std_logic_vector (3 downto 0);
        card1_5 : in std_logic_vector (3 downto 0);
        money1  : in std_logic_vector (10 downto 0);
	split1 	: in std_logic;
	bet1 : in std_logic_vector (1 downto 0);
	doubledown1 : in std_logic;
	insurance1	: in std_logic;

        player_b : in std_logic;
        card2_1 : in std_logic_vector (3 downto 0);
        card2_2 : in std_logic_vector (3 downto 0);
        card2_3 : in std_logic_vector (3 downto 0);
        card2_4 : in std_logic_vector (3 downto 0);
        card2_5 : in std_logic_vector (3 downto 0);
        money2  : in std_logic_vector (10 downto 0);
	split2	: in std_logic;
bet2 : in std_logic_vector (1 downto 0);
	doubledown2 : in std_logic;
	insurance2	: in std_logic;

        player_c : in std_logic;
        card3_1 : in std_logic_vector (3 downto 0);
        card3_2 : in std_logic_vector (3 downto 0);
        card3_3 : in std_logic_vector (3 downto 0);
        card3_4 : in std_logic_vector (3 downto 0);
        card3_5 : in std_logic_vector (3 downto 0);
        money3  : in std_logic_vector (10 downto 0);
	split3	: in std_logic;
	bet3 : in std_logic_vector (1 downto 0);
	doubledown3 : in std_logic;
	insurance3	: in std_logic;

        player_d : in std_logic;
        card4_1 : in std_logic_vector (3 downto 0);
        card4_2 : in std_logic_vector (3 downto 0);
        card4_3 : in std_logic_vector (3 downto 0);
        card4_4 : in std_logic_vector (3 downto 0);
        card4_5 : in std_logic_vector (3 downto 0);
        money4  : in std_logic_vector (10 downto 0);
	split4	: in std_logic;
	bet4 : in std_logic_vector (1 downto 0);
	doubledown4 : in std_logic;
	insurance4	: in std_logic;
	        card5_1 : in std_logic_vector (3 downto 0);
        card5_2 : in std_logic_vector (3 downto 0);
        card5_3 : in std_logic_vector (3 downto 0);
        card5_4 : in std_logic_vector (3 downto 0);
        card5_5 : in std_logic_vector (3 downto 0);
		  split1_1: in std_logic_vector (3 downto 0);
		  split1_2: in std_logic_vector (3 downto 0);
		  split1_3 : in std_logic_vector (3 downto 0);
		  split1_4: in std_logic_vector (3 downto 0);
		  split1_5: in std_logic_vector (3 downto 0);
		  
split2_1: in std_logic_vector (3 downto 0);
 split2_2: in std_logic_vector (3 downto 0);
 split2_3: in std_logic_vector (3 downto 0);
 split2_4: in std_logic_vector (3 downto 0);
 split2_5: in std_logic_vector (3 downto 0);
 split3_1: in std_logic_vector (3 downto 0);
 split3_2: in std_logic_vector (3 downto 0);
 split3_3: in std_logic_vector (3 downto 0);
 split3_4: in std_logic_vector (3 downto 0);
 split3_5: in std_logic_vector (3 downto 0);
 split4_1: in std_logic_vector (3 downto 0);
 split4_2: in std_logic_vector (3 downto 0);
 split4_3: in std_logic_vector (3 downto 0);
 split4_4: in std_logic_vector (3 downto 0);
 split4_5 : in std_logic_vector (3 downto 0)
);
end main;

