djkahgydubauid
