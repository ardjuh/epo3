entity gpu_driver_tb is
end entity;