library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of graphics_driver_tb is
component graphics_driver
	 port (
        h_pos : in std_logic_vector(9 downto 0);
        v_pos : in std_logic_vector(9 downto 0);
        red   : out std_logic_vector(3 downto 0);
        green : out std_logic_vector(3 downto 0);
        blue  : out std_logic_vector(3 downto 0));
end component;

signal h_pos: std_logic_vector(9 downto 0);
signal v_pos: std_logic_vector(9 downto 0);
signal red: std_logic_vector(3 downto 0);
signal green: std_logic_vector(3 downto 0);
signal blue: std_logic_vector(3 downto 0);


begin
test: graphics_driver port map (h_pos,v_pos,red,green,blue);

h_pos <= "0000000000" after 0 ns,
"0000000001" after 40 ns,
"0000000010" after 80 ns,
"0000000011" after 120 ns,
"0000000100" after 160 ns,
"0000000101" after 200 ns,
"0000000110" after 240 ns,
"0000000111" after 280 ns,
"0000001000" after 320 ns,
"0000001001" after 360 ns,
"0000001010" after 400 ns,
"0000001011" after 440 ns,
"0000001100" after 480 ns,
"0000001101" after 520 ns,
"0000001110" after 560 ns,
"0000001111" after 600 ns,
"0000010000" after 640 ns,
"0000010001" after 680 ns,
"0000010010" after 720 ns,
"0000010011" after 760 ns,
"0000010100" after 800 ns,
"0000010101" after 840 ns,
"0000010110" after 880 ns,
"0000010111" after 920 ns,
"0000011000" after 960 ns,
"0000011001" after 1000 ns,
"0000011010" after 1040 ns,
"0000011011" after 1080 ns,
"0000011100" after 1120 ns,
"0000011101" after 1160 ns,
"0000011110" after 1200 ns,
"0000011111" after 1240 ns,
"0000100000" after 1280 ns,
"0000100001" after 1320 ns,
"0000100010" after 1360 ns,
"0000100011" after 1400 ns,
"0000100100" after 1440 ns,
"0000100101" after 1480 ns,
"0000100110" after 1520 ns,
"0000100111" after 1560 ns,
"0000101000" after 1600 ns,
"0000101001" after 1640 ns,
"0000101010" after 1680 ns,
"0000101011" after 1720 ns,
"0000101100" after 1760 ns,
"0000101101" after 1800 ns,
"0000101110" after 1840 ns,
"0000101111" after 1880 ns,
"0000110000" after 1920 ns,
"0000110001" after 1960 ns,
"0000110010" after 2000 ns,
"0000110011" after 2040 ns,
"0000110100" after 2080 ns,
"0000110101" after 2120 ns,
"0000110110" after 2160 ns,
"0000110111" after 2200 ns,
"0000111000" after 2240 ns,
"0000111001" after 2280 ns,
"0000111010" after 2320 ns,
"0000111011" after 2360 ns,
"0000111100" after 2400 ns,
"0000111101" after 2440 ns,
"0000111110" after 2480 ns,
"0000111111" after 2520 ns,
"0001000000" after 2560 ns,
"0001000001" after 2600 ns,
"0001000010" after 2640 ns,
"0001000011" after 2680 ns,
"0001000100" after 2720 ns,
"0001000101" after 2760 ns,
"0001000110" after 2800 ns,
"0001000111" after 2840 ns,
"0001001000" after 2880 ns,
"0001001001" after 2920 ns,
"0001001010" after 2960 ns,
"0001001011" after 3000 ns,
"0001001100" after 3040 ns,
"0001001101" after 3080 ns,
"0001001110" after 3120 ns,
"0001001111" after 3160 ns,
"0001010000" after 3200 ns,
"0001010001" after 3240 ns,
"0001010010" after 3280 ns,
"0001010011" after 3320 ns,
"0001010100" after 3360 ns,
"0001010101" after 3400 ns,
"0001010110" after 3440 ns,
"0001010111" after 3480 ns,
"0001011000" after 3520 ns,
"0001011001" after 3560 ns,
"0001011010" after 3600 ns,
"0001011011" after 3640 ns,
"0001011100" after 3680 ns,
"0001011101" after 3720 ns,
"0001011110" after 3760 ns,
"0001011111" after 3800 ns,
"0001100000" after 3840 ns,
"0001100001" after 3880 ns,
"0001100010" after 3920 ns,
"0001100011" after 3960 ns,
"0001100100" after 4000 ns,
"0001100101" after 4040 ns,
"0001100110" after 4080 ns,
"0001100111" after 4120 ns,
"0001101000" after 4160 ns,
"0001101001" after 4200 ns,
"0001101010" after 4240 ns,
"0001101011" after 4280 ns,
"0001101100" after 4320 ns,
"0001101101" after 4360 ns,
"0001101110" after 4400 ns,
"0001101111" after 4440 ns,
"0001110000" after 4480 ns,
"0001110001" after 4520 ns,
"0001110010" after 4560 ns,
"0001110011" after 4600 ns,
"0001110100" after 4640 ns,
"0001110101" after 4680 ns,
"0001110110" after 4720 ns,
"0001110111" after 4760 ns,
"0001111000" after 4800 ns,
"0001111001" after 4840 ns,
"0001111010" after 4880 ns,
"0001111011" after 4920 ns,
"0001111100" after 4960 ns,
"0001111101" after 5000 ns,
"0001111110" after 5040 ns,
"0001111111" after 5080 ns,
"0010000000" after 5120 ns,
"0010000001" after 5160 ns,
"0010000010" after 5200 ns,
"0010000011" after 5240 ns,
"0010000100" after 5280 ns,
"0010000101" after 5320 ns,
"0010000110" after 5360 ns,
"0010000111" after 5400 ns,
"0010001000" after 5440 ns,
"0010001001" after 5480 ns,
"0010001010" after 5520 ns,
"0010001011" after 5560 ns,
"0010001100" after 5600 ns,
"0010001101" after 5640 ns,
"0010001110" after 5680 ns,
"0010001111" after 5720 ns,
"0010010000" after 5760 ns,
"0010010001" after 5800 ns,
"0010010010" after 5840 ns,
"0010010011" after 5880 ns,
"0010010100" after 5920 ns,
"0010010101" after 5960 ns,
"0010010110" after 6000 ns,
"0010010111" after 6040 ns,
"0010011000" after 6080 ns,
"0010011001" after 6120 ns,
"0010011010" after 6160 ns,
"0010011011" after 6200 ns,
"0010011100" after 6240 ns,
"0010011101" after 6280 ns,
"0010011110" after 6320 ns,
"0010011111" after 6360 ns,
"0010100000" after 6400 ns,
"0010100001" after 6440 ns,
"0010100010" after 6480 ns,
"0010100011" after 6520 ns,
"0010100100" after 6560 ns,
"0010100101" after 6600 ns,
"0010100110" after 6640 ns,
"0010100111" after 6680 ns,
"0010101000" after 6720 ns,
"0010101001" after 6760 ns,
"0010101010" after 6800 ns,
"0010101011" after 6840 ns,
"0010101100" after 6880 ns,
"0010101101" after 6920 ns,
"0010101110" after 6960 ns,
"0010101111" after 7000 ns,
"0010110000" after 7040 ns,
"0010110001" after 7080 ns,
"0010110010" after 7120 ns,
"0010110011" after 7160 ns,
"0010110100" after 7200 ns,
"0010110101" after 7240 ns,
"0010110110" after 7280 ns,
"0010110111" after 7320 ns,
"0010111000" after 7360 ns,
"0010111001" after 7400 ns,
"0010111010" after 7440 ns,
"0010111011" after 7480 ns,
"0010111100" after 7520 ns,
"0010111101" after 7560 ns,
"0010111110" after 7600 ns,
"0010111111" after 7640 ns,
"0011000000" after 7680 ns,
"0011000001" after 7720 ns,
"0011000010" after 7760 ns,
"0011000011" after 7800 ns,
"0011000100" after 7840 ns,
"0011000101" after 7880 ns,
"0011000110" after 7920 ns,
"0011000111" after 7960 ns,
"0011001000" after 8000 ns,
"0011001001" after 8040 ns,
"0011001010" after 8080 ns,
"0011001011" after 8120 ns,
"0011001100" after 8160 ns,
"0011001101" after 8200 ns,
"0011001110" after 8240 ns,
"0011001111" after 8280 ns,
"0011010000" after 8320 ns,
"0011010001" after 8360 ns,
"0011010010" after 8400 ns,
"0011010011" after 8440 ns,
"0011010100" after 8480 ns,
"0011010101" after 8520 ns,
"0011010110" after 8560 ns,
"0011010111" after 8600 ns,
"0011011000" after 8640 ns,
"0011011001" after 8680 ns,
"0011011010" after 8720 ns,
"0011011011" after 8760 ns,
"0011011100" after 8800 ns,
"0011011101" after 8840 ns,
"0011011110" after 8880 ns,
"0011011111" after 8920 ns,
"0011100000" after 8960 ns,
"0011100001" after 9000 ns,
"0011100010" after 9040 ns,
"0011100011" after 9080 ns,
"0011100100" after 9120 ns,
"0011100101" after 9160 ns,
"0011100110" after 9200 ns,
"0011100111" after 9240 ns,
"0011101000" after 9280 ns,
"0011101001" after 9320 ns,
"0011101010" after 9360 ns,
"0011101011" after 9400 ns,
"0011101100" after 9440 ns,
"0011101101" after 9480 ns,
"0011101110" after 9520 ns,
"0011101111" after 9560 ns,
"0011110000" after 9600 ns,
"0011110001" after 9640 ns,
"0011110010" after 9680 ns,
"0011110011" after 9720 ns,
"0011110100" after 9760 ns,
"0011110101" after 9800 ns,
"0011110110" after 9840 ns,
"0011110111" after 9880 ns,
"0011111000" after 9920 ns,
"0011111001" after 9960 ns,
"0011111010" after 10000 ns,
"0011111011" after 10040 ns,
"0011111100" after 10080 ns,
"0011111101" after 10120 ns,
"0011111110" after 10160 ns,
"0011111111" after 10200 ns,
"0100000000" after 10240 ns,
"0100000001" after 10280 ns,
"0100000010" after 10320 ns,
"0100000011" after 10360 ns,
"0100000100" after 10400 ns,
"0100000101" after 10440 ns,
"0100000110" after 10480 ns,
"0100000111" after 10520 ns,
"0100001000" after 10560 ns,
"0100001001" after 10600 ns,
"0100001010" after 10640 ns,
"0100001011" after 10680 ns,
"0100001100" after 10720 ns,
"0100001101" after 10760 ns,
"0100001110" after 10800 ns,
"0100001111" after 10840 ns,
"0100010000" after 10880 ns,
"0100010001" after 10920 ns,
"0100010010" after 10960 ns,
"0100010011" after 11000 ns,
"0100010100" after 11040 ns,
"0100010101" after 11080 ns,
"0100010110" after 11120 ns,
"0100010111" after 11160 ns,
"0100011000" after 11200 ns,
"0100011001" after 11240 ns,
"0100011010" after 11280 ns,
"0100011011" after 11320 ns,
"0100011100" after 11360 ns,
"0100011101" after 11400 ns,
"0100011110" after 11440 ns,
"0100011111" after 11480 ns,
"0100100000" after 11520 ns,
"0100100001" after 11560 ns,
"0100100010" after 11600 ns,
"0100100011" after 11640 ns,
"0100100100" after 11680 ns,
"0100100101" after 11720 ns,
"0100100110" after 11760 ns,
"0100100111" after 11800 ns,
"0100101000" after 11840 ns,
"0100101001" after 11880 ns,
"0100101010" after 11920 ns,
"0100101011" after 11960 ns,
"0100101100" after 12000 ns,
"0100101101" after 12040 ns,
"0100101110" after 12080 ns,
"0100101111" after 12120 ns,
"0100110000" after 12160 ns,
"0100110001" after 12200 ns,
"0100110010" after 12240 ns,
"0100110011" after 12280 ns,
"0100110100" after 12320 ns,
"0100110101" after 12360 ns,
"0100110110" after 12400 ns,
"0100110111" after 12440 ns,
"0100111000" after 12480 ns,
"0100111001" after 12520 ns,
"0100111010" after 12560 ns,
"0100111011" after 12600 ns,
"0100111100" after 12640 ns,
"0100111101" after 12680 ns,
"0100111110" after 12720 ns,
"0100111111" after 12760 ns,
"0101000000" after 12800 ns,
"0101000001" after 12840 ns,
"0101000010" after 12880 ns,
"0101000011" after 12920 ns,
"0101000100" after 12960 ns,
"0101000101" after 13000 ns,
"0101000110" after 13040 ns,
"0101000111" after 13080 ns,
"0101001000" after 13120 ns,
"0101001001" after 13160 ns,
"0101001010" after 13200 ns,
"0101001011" after 13240 ns,
"0101001100" after 13280 ns,
"0101001101" after 13320 ns,
"0101001110" after 13360 ns,
"0101001111" after 13400 ns,
"0101010000" after 13440 ns,
"0101010001" after 13480 ns,
"0101010010" after 13520 ns,
"0101010011" after 13560 ns,
"0101010100" after 13600 ns,
"0101010101" after 13640 ns,
"0101010110" after 13680 ns,
"0101010111" after 13720 ns,
"0101011000" after 13760 ns,
"0101011001" after 13800 ns,
"0101011010" after 13840 ns,
"0101011011" after 13880 ns,
"0101011100" after 13920 ns,
"0101011101" after 13960 ns,
"0101011110" after 14000 ns,
"0101011111" after 14040 ns,
"0101100000" after 14080 ns,
"0101100001" after 14120 ns,
"0101100010" after 14160 ns,
"0101100011" after 14200 ns,
"0101100100" after 14240 ns,
"0101100101" after 14280 ns,
"0101100110" after 14320 ns,
"0101100111" after 14360 ns,
"0101101000" after 14400 ns,
"0101101001" after 14440 ns,
"0101101010" after 14480 ns,
"0101101011" after 14520 ns,
"0101101100" after 14560 ns,
"0101101101" after 14600 ns,
"0101101110" after 14640 ns,
"0101101111" after 14680 ns,
"0101110000" after 14720 ns,
"0101110001" after 14760 ns,
"0101110010" after 14800 ns,
"0101110011" after 14840 ns,
"0101110100" after 14880 ns,
"0101110101" after 14920 ns,
"0101110110" after 14960 ns,
"0101110111" after 15000 ns,
"0101111000" after 15040 ns,
"0101111001" after 15080 ns,
"0101111010" after 15120 ns,
"0101111011" after 15160 ns,
"0101111100" after 15200 ns,
"0101111101" after 15240 ns,
"0101111110" after 15280 ns,
"0101111111" after 15320 ns,
"0110000000" after 15360 ns,
"0110000001" after 15400 ns,
"0110000010" after 15440 ns,
"0110000011" after 15480 ns,
"0110000100" after 15520 ns,
"0110000101" after 15560 ns,
"0110000110" after 15600 ns,
"0110000111" after 15640 ns,
"0110001000" after 15680 ns,
"0110001001" after 15720 ns,
"0110001010" after 15760 ns,
"0110001011" after 15800 ns,
"0110001100" after 15840 ns,
"0110001101" after 15880 ns,
"0110001110" after 15920 ns,
"0110001111" after 15960 ns,
"0110010000" after 16000 ns,
"0110010001" after 16040 ns,
"0110010010" after 16080 ns,
"0110010011" after 16120 ns,
"0110010100" after 16160 ns,
"0110010101" after 16200 ns,
"0110010110" after 16240 ns,
"0110010111" after 16280 ns,
"0110011000" after 16320 ns,
"0110011001" after 16360 ns,
"0110011010" after 16400 ns,
"0110011011" after 16440 ns,
"0110011100" after 16480 ns,
"0110011101" after 16520 ns,
"0110011110" after 16560 ns,
"0110011111" after 16600 ns,
"0110100000" after 16640 ns,
"0110100001" after 16680 ns,
"0110100010" after 16720 ns,
"0110100011" after 16760 ns,
"0110100100" after 16800 ns,
"0110100101" after 16840 ns,
"0110100110" after 16880 ns,
"0110100111" after 16920 ns,
"0110101000" after 16960 ns,
"0110101001" after 17000 ns,
"0110101010" after 17040 ns,
"0110101011" after 17080 ns,
"0110101100" after 17120 ns,
"0110101101" after 17160 ns,
"0110101110" after 17200 ns,
"0110101111" after 17240 ns,
"0110110000" after 17280 ns,
"0110110001" after 17320 ns,
"0110110010" after 17360 ns,
"0110110011" after 17400 ns,
"0110110100" after 17440 ns,
"0110110101" after 17480 ns,
"0110110110" after 17520 ns,
"0110110111" after 17560 ns,
"0110111000" after 17600 ns,
"0110111001" after 17640 ns,
"0110111010" after 17680 ns,
"0110111011" after 17720 ns,
"0110111100" after 17760 ns,
"0110111101" after 17800 ns,
"0110111110" after 17840 ns,
"0110111111" after 17880 ns,
"0111000000" after 17920 ns,
"0111000001" after 17960 ns,
"0111000010" after 18000 ns,
"0111000011" after 18040 ns,
"0111000100" after 18080 ns,
"0111000101" after 18120 ns,
"0111000110" after 18160 ns,
"0111000111" after 18200 ns,
"0111001000" after 18240 ns,
"0111001001" after 18280 ns,
"0111001010" after 18320 ns,
"0111001011" after 18360 ns,
"0111001100" after 18400 ns,
"0111001101" after 18440 ns,
"0111001110" after 18480 ns,
"0111001111" after 18520 ns,
"0111010000" after 18560 ns,
"0111010001" after 18600 ns,
"0111010010" after 18640 ns,
"0111010011" after 18680 ns,
"0111010100" after 18720 ns,
"0111010101" after 18760 ns,
"0111010110" after 18800 ns,
"0111010111" after 18840 ns,
"0111011000" after 18880 ns,
"0111011001" after 18920 ns,
"0111011010" after 18960 ns,
"0111011011" after 19000 ns,
"0111011100" after 19040 ns,
"0111011101" after 19080 ns,
"0111011110" after 19120 ns,
"0111011111" after 19160 ns,
"0111100000" after 19200 ns,
"0111100001" after 19240 ns,
"0111100010" after 19280 ns,
"0111100011" after 19320 ns,
"0111100100" after 19360 ns,
"0111100101" after 19400 ns,
"0111100110" after 19440 ns,
"0111100111" after 19480 ns,
"0111101000" after 19520 ns,
"0111101001" after 19560 ns,
"0111101010" after 19600 ns,
"0111101011" after 19640 ns,
"0111101100" after 19680 ns,
"0111101101" after 19720 ns,
"0111101110" after 19760 ns,
"0111101111" after 19800 ns,
"0111110000" after 19840 ns,
"0111110001" after 19880 ns,
"0111110010" after 19920 ns,
"0111110011" after 19960 ns,
"0111110100" after 20000 ns,
"0111110101" after 20040 ns,
"0111110110" after 20080 ns,
"0111110111" after 20120 ns,
"0111111000" after 20160 ns,
"0111111001" after 20200 ns,
"0111111010" after 20240 ns,
"0111111011" after 20280 ns,
"0111111100" after 20320 ns,
"0111111101" after 20360 ns,
"0111111110" after 20400 ns,
"0111111111" after 20440 ns,
"1000000000" after 20480 ns,
"1000000001" after 20520 ns,
"1000000010" after 20560 ns,
"1000000011" after 20600 ns,
"1000000100" after 20640 ns,
"1000000101" after 20680 ns,
"1000000110" after 20720 ns,
"1000000111" after 20760 ns,
"1000001000" after 20800 ns,
"1000001001" after 20840 ns,
"1000001010" after 20880 ns,
"1000001011" after 20920 ns,
"1000001100" after 20960 ns,
"1000001101" after 21000 ns,
"1000001110" after 21040 ns,
"1000001111" after 21080 ns,
"1000010000" after 21120 ns,
"1000010001" after 21160 ns,
"1000010010" after 21200 ns,
"1000010011" after 21240 ns,
"1000010100" after 21280 ns,
"1000010101" after 21320 ns,
"1000010110" after 21360 ns,
"1000010111" after 21400 ns,
"1000011000" after 21440 ns,
"1000011001" after 21480 ns,
"1000011010" after 21520 ns,
"1000011011" after 21560 ns,
"1000011100" after 21600 ns,
"1000011101" after 21640 ns,
"1000011110" after 21680 ns,
"1000011111" after 21720 ns,
"1000100000" after 21760 ns,
"1000100001" after 21800 ns,
"1000100010" after 21840 ns,
"1000100011" after 21880 ns,
"1000100100" after 21920 ns,
"1000100101" after 21960 ns,
"1000100110" after 22000 ns,
"1000100111" after 22040 ns,
"1000101000" after 22080 ns,
"1000101001" after 22120 ns,
"1000101010" after 22160 ns,
"1000101011" after 22200 ns,
"1000101100" after 22240 ns,
"1000101101" after 22280 ns,
"1000101110" after 22320 ns,
"1000101111" after 22360 ns,
"1000110000" after 22400 ns,
"1000110001" after 22440 ns,
"1000110010" after 22480 ns,
"1000110011" after 22520 ns,
"1000110100" after 22560 ns,
"1000110101" after 22600 ns,
"1000110110" after 22640 ns,
"1000110111" after 22680 ns,
"1000111000" after 22720 ns,
"1000111001" after 22760 ns,
"1000111010" after 22800 ns,
"1000111011" after 22840 ns,
"1000111100" after 22880 ns,
"1000111101" after 22920 ns,
"1000111110" after 22960 ns,
"1000111111" after 23000 ns,
"1001000000" after 23040 ns,
"1001000001" after 23080 ns,
"1001000010" after 23120 ns,
"1001000011" after 23160 ns,
"1001000100" after 23200 ns,
"1001000101" after 23240 ns,
"1001000110" after 23280 ns,
"1001000111" after 23320 ns,
"1001001000" after 23360 ns,
"1001001001" after 23400 ns,
"1001001010" after 23440 ns,
"1001001011" after 23480 ns,
"1001001100" after 23520 ns,
"1001001101" after 23560 ns,
"1001001110" after 23600 ns,
"1001001111" after 23640 ns,
"1001010000" after 23680 ns,
"1001010001" after 23720 ns,
"1001010010" after 23760 ns,
"1001010011" after 23800 ns,
"1001010100" after 23840 ns,
"1001010101" after 23880 ns,
"1001010110" after 23920 ns,
"1001010111" after 23960 ns,
"1001011000" after 24000 ns,
"1001011001" after 24040 ns,
"1001011010" after 24080 ns,
"1001011011" after 24120 ns,
"1001011100" after 24160 ns,
"1001011101" after 24200 ns,
"1001011110" after 24240 ns,
"1001011111" after 24280 ns,
"1001100000" after 24320 ns,
"1001100001" after 24360 ns,
"1001100010" after 24400 ns,
"1001100011" after 24440 ns,
"1001100100" after 24480 ns,
"1001100101" after 24520 ns,
"1001100110" after 24560 ns,
"1001100111" after 24600 ns,
"1001101000" after 24640 ns,
"1001101001" after 24680 ns,
"1001101010" after 24720 ns,
"1001101011" after 24760 ns,
"1001101100" after 24800 ns,
"1001101101" after 24840 ns,
"1001101110" after 24880 ns,
"1001101111" after 24920 ns,
"1001110000" after 24960 ns,
"1001110001" after 25000 ns,
"1001110010" after 25040 ns,
"1001110011" after 25080 ns,
"1001110100" after 25120 ns,
"1001110101" after 25160 ns,
"1001110110" after 25200 ns,
"1001110111" after 25240 ns,
"1001111000" after 25280 ns,
"1001111001" after 25320 ns,
"1001111010" after 25360 ns,
"1001111011" after 25400 ns,
"1001111100" after 25440 ns,
"1001111101" after 25480 ns,
"1001111110" after 25520 ns,
"1001111111" after 25560 ns;

end behaviour;
