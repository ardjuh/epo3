library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


entity counter is
	port(
	clk: in std_logic;
	reset: in std_logic;
	x_pos: out std_logic_vector(9 downto 0);
	y_pos: out std_logic_vector(9 downto 0));
end counter;

